library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity control_unit is
  port (
  );
end entity;

architecture behave of control_unit is
begin
end architecture;

